** Profile: "SCHEMATIC1-test1234"  [ c:\users\skypv\desktop\p1_2025_433d_dinca_matei_gsd_tema_11_orcad\p1_2025_433d_dinca_matei_gsd_tema_11_orcad\schematics\test123-pspicefiles\schematic1\test1234.sim ] 

** Creating circuit file "test1234.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../MovedFiles/bc846b.lib" 
.LIB "../../../MovedFiles/bc856b.lib" 
* From [PSPICE NETLIST] section of C:\Users\skypv\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 2ms 0 1u SKIPBP 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
